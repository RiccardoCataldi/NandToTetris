module alu(input [15:0] x, input [15:0] y, input zx,input nx,input zy,input ny,input f,input no,output [15:0] out, output zr,output ng);
endmodule
