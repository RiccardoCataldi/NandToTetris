module not16(input [15:0] in, output [15:0] out);
    not2 n0(.a(in[0]), .y(out[0]));
    not2 n1(.a(in[1]), .y(out[1]));
    not2 n2(.a(in[2]), .y(out[2]));
    not2 n3(.a(in[3]), .y(out[3]));
    not2 n4(.a(in[4]), .y(out[4]));
    not2 n5(.a(in[5]), .y(out[5]));
    not2 n6(.a(in[6]), .y(out[6]));
    not2 n7(.a(in[7]), .y(out[7]));
    not2 n8(.a(in[8]), .y(out[8]));
    not2 n9(.a(in[9]), .y(out[9]));
    not2 n10(.a(in[10]), .y(out[10]));
    not2 n11(.a(in[11]), .y(out[11]));
    not2 n12(.a(in[12]), .y(out[12]));
    not2 n13(.a(in[13]), .y(out[13]));
    not2 n14(.a(in[14]), .y(out[14]));
    not2 n15(.a(in[15]), .y(out[15]));
endmodule
